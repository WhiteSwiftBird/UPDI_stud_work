//////////////////////////////////////////////////////////////////////////////////
// Company: POLYTHEC
// Engineer: ARTEM
// 
// Create Date: 25.06.2025 00:17:38
// Design Name: UPDI Physical level
// Module Name: PHY
// Project Name: 
// Target Devices: UPDI
// Tool Versions: 
// Description: PHY level of UPDI, w/r info in AVR
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module PHY (

	input clk,
	input rst,
	input ten, //transmission enable
	input ren,
	output csb0,
	output web0,
	output [6:0]  addr0,
	inout logic [11:0] io_data,
	output tend,  //end-transmission signal
	output rend  //end-receiving signal
	
	);
	
	logic pwdata, prdata;
	
	PHY_LOADER loader_from_mem ( 
	
	                             .clk(clk),
										  .rst(rst), 
	                             .ten(ten), 
										  .ren(ren), 
										  .csb0(csb0), 
										  .web0(web0), 
										  .addr0(addr0), 
										  .io_data(io_data), 
										  .pwdata(pwdata), 
										  .prdata(prdata),
										  .tend(tend),
										  .rend(rend) 
										  
										);
	
	/*apb_uart UART              ( 
	
	                             .pwdata(pwdata), 
	                             .prdata(prdata) 
										  
										);*/
										
endmodule
										
module top_UPDI (

);
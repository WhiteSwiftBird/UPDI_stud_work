//////////////////////////////////////////////////////////////////////////////////
// Company: POLYTHEC
// Engineer: ARTEM
// 
// Create Date: 26.06.2025 00:17:38
// Design Name: PHY rx testbench 
// Module Name: PHY_tb_rx
// Project Name: 
// Target Devices: UPDI
// Tool Versions: 
// Description: testbench of PHY level receiving of UPDI
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: Пока не подключен полноценный UART внутренние сигналы PHY нужно выводить наружу для проверки правильности отправки данных
// 
//////////////////////////////////////////////////////////////////////////////////

`timescale 10ps / 1ps

module PHY_tb_rx ;

    logic clk;
    logic rst;
    logic ten; 
    logic ren;
    logic csb0;
    logic web0;
    logic [6:0]  addr0;
    logic [11:0] i_data;
    logic [11:0] o_data;	 
    logic tend; 
    logic rend;  
    logic pwdata; 
    logic prdata; 
	
    int iterator, error, cnt, one_delay; //variables cnt is a immitation of getting data from mem
	 
	 logic [2:0] tv [1000:0]; //testvector
    logic [11:0] o_data_reg;
    PHY_LOADER uut (
               .clk(clk),
               .rst(rst), 
               .ten(ten), 
               .ren(ren), 
               .csb0(csb0), 
               .web0(web0), 
               .addr0(addr0), 
					.i_data(i_data),
					.o_data(o_data), 
               .pwdata(pwdata), 
               .prdata(prdata),
               .tend(tend),
               .rend(rend) 
            );
				
				
				
				
    initial 
      begin
		  
		  //variables init
		  $readmemb("D:/UPDI Project RADAR/UPDI_stud_work/src/PHY/PHY_tb_rx.tv", tv);
		  iterator = 0;
		  cnt = 0;
		  error = 0;
		  one_delay = 0;
		  
		  //uut signals init
		  { ten, ren, prdata } = tv [0];
		  //rst = 0;
		  clk = 1;
		  //#5;
		  //rst = 1;
		  
      end
		
		
    always 
      begin
		  
        #5;
        clk = ~clk;
		
      end
		
		
    always @(posedge clk)
      begin
				
				o_data_reg[(cnt % 12)] <= prdata;
				
				if (one_delay > 0)
				cnt <= cnt + 1; 
				
				one_delay += 1;
			 
			 
		  if ( tv [cnt] === 'x )
		    begin
				
				  $display ("Test ended in %d iterations and handle %d errors", cnt + 1, error);
				  $stop;
				  
			 end
	     
	   end
		
    always @(negedge clk)
	 
	   begin
	 
	       { ten, ren, prdata } <= tv [cnt];
			 
		    if (cnt % 12 == 0)
		    begin
			 
			   if ( o_data != o_data_reg)
			 
			       begin
				
				    $error ("Error detected in %d line", iterator);
				    error += 1;
				    iterator += 1;
				
				    end
				
			 end
			 
		end
		
		
endmodule
1_0_101000101010
1_0_111100001111
1_0_010100101000
1_0_100000000001
1_0_111101000110
//////////////////////////////////////////////////////////////////////////////////
// Company: POLYTHEC
// Engineer: ARTEM
// 
// Create Date: 25.06.2025 00:17:38
// Design Name: UPDI Physical level loader
// Module Name: PHY_LOADER
// Project Name: 
// Target Devices: UPDI
// Tool Versions: 
// Description: Loader of prepared in CG data, use UART to t/r data to AVR
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module PHY_LOADER (
	
     input clk,
	  input rst,   //reset while start UPDI
     input logic ten,  //transmission enable
     input logic ren, //receive enable
	 //input ACK, //acknowledge bit, unnecessary
    output logic csb0,
    output logic web0,
    output logic [6:0]  addr0,
	  input logic [11:0] i_data,
	 output logic [11:0] o_data, //не забыть положить сюда данные, в самом топовом модуле соединить соответсвующий выход с память BUFF_MEM
	  input logic prdata, //RX UART
	 output logic pwdata,  //TX UART
	 output logic tend,  //end-transmission signal
	 output logic rend  //end-receiving signal	 
	
    );
	
	logic [11:0] io_data_reg;
	logic [3:0]  counter;
	
	enum logic [1:0] {IDLE = 2'b00, TR = 2'b01, RC = 2'b10} state, next_state;
	
	
	
	always_ff @(posedge clk)
	  if (!rst)
	    state <= IDLE;
	  else
	    state <= next_state;
	
	
   always_comb
	  begin
		
		 next_state = state;
		
		 case (state)
		    
			 IDLE:      if (!ten)
			            next_state = TR;
						  
					      else if (!ren)
					      next_state = RC;
						  
			 TR:        if (!tend && !ren)
			            next_state = RC;
							
						   else if (!tend && ren)
						   next_state = IDLE;
						  
			 RC:        if (!rend)
			            next_state = IDLE;
						  
			 default:   next_state = IDLE;
		
		 endcase 
		
	  end
	
   always_ff @(negedge clk)
      begin
		  
		  case (state)
		  
            IDLE: begin
				
				        csb0 <= 1'b1;
				        counter <= '0;
						  addr0 <= '0;
						  tend <= 1'b0;
						  rend <= 1'b0;
		              io_data_reg <= '0;
						  
			         end
			   //transmission
            TR:   begin
				        if (counter == 0)
						    begin
							 
							   csb0 <= 1'b0;
							   web0 <= 1'b1;
						      //io_data_reg [11:0] <= i_data [11:0];
								
							 end
						  
	                 if (counter < 12)
				          begin
				
				            pwdata <= i_data[counter];
					         //i_data <= (i_data >> 1);
					         counter <= counter + 1;
					 
					       end
					 
				        else
				          begin
					  
					         counter <= '0;
                        addr0 <= addr0 + 1;
					  
					       end
					  
				        //end of transmission
				        if ( (&addr0) && (counter == 12) )
				          begin 
					  
					         addr0 <= '0;
					         tend <= 1'b0;
					  
					       end
				        else
				            tend <= 1'b1;	
					
			
	               end 
						
				//receiving	
            RC:   begin
				        if (counter < 12)
						    begin
							 
							   io_data_reg [counter] <= prdata;
								counter <= counter + 1;
								
							 end
							 
				        else
				          begin
					         
								csb0 <= 1'b0;
								web0 <= 1'b0;
								o_data <= io_data_reg;
					         counter <= 1'b0;
                        addr0 <= addr0 + 1;
					  
					       end
							 
				        if ( (&addr0) && (counter == 11) )
				          begin 
					  
					         addr0 <= '0;
					         rend <= 1'b0;
					  
					       end
				        else
				            rend <= 1'b1;	
						  
						  
						end
				
            default: begin
				
				           csb0 = 1'b1;
				           counter = '0;
						     addr0 = '0;
						     tend = 1'b0;
						     rend = 1'b0;
		                 io_data_reg = '0;
							  
			            end
			endcase
		
		  
        end
			     
		  
endmodule